module RAM(in, address, load, out);
